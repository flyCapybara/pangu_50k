module moduleName (
    input wire a,
    input wire b,
    output wire y
);
    
endmodule